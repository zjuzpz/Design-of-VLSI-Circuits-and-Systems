module NLC_32ch (
input [31:0] ch0_coeff_1_0,
input [31:0] ch0_coeff_1_1,
input [31:0] ch0_coeff_1_2,
input [31:0] ch0_coeff_1_3,
input [31:0] ch0_coeff_1_4,
input [31:0] ch0_coeff_1_5,
input [31:0] ch0_coeff_1_6,
input [31:0] ch0_coeff_1_7,
input [31:0] ch0_coeff_1_8,
input [31:0] ch0_coeff_1_9,
input [31:0] ch0_coeff_1_10,
input [31:0] ch0_coeff_2_0,
input [31:0] ch0_coeff_2_1,
input [31:0] ch0_coeff_2_2,
input [31:0] ch0_coeff_2_3,
input [31:0] ch0_coeff_2_4,
input [31:0] ch0_coeff_2_5,
input [31:0] ch0_coeff_2_6,
input [31:0] ch0_coeff_2_7,
input [31:0] ch0_coeff_2_8,
input [31:0] ch0_coeff_2_9,
input [31:0] ch0_coeff_2_10,
input [31:0] ch0_coeff_3_0,
input [31:0] ch0_coeff_3_1,
input [31:0] ch0_coeff_3_2,
input [31:0] ch0_coeff_3_3,
input [31:0] ch0_coeff_3_4,
input [31:0] ch0_coeff_3_5,
input [31:0] ch0_coeff_3_6,
input [31:0] ch0_coeff_3_7,
input [31:0] ch0_coeff_3_8,
input [31:0] ch0_coeff_3_9,
input [31:0] ch0_coeff_3_10,
input [31:0] ch0_coeff_4_0,
input [31:0] ch0_coeff_4_1,
input [31:0] ch0_coeff_4_2,
input [31:0] ch0_coeff_4_3,
input [31:0] ch0_coeff_4_4,
input [31:0] ch0_coeff_4_5,
input [31:0] ch0_coeff_4_6,
input [31:0] ch0_coeff_4_7,
input [31:0] ch0_coeff_4_8,
input [31:0] ch0_coeff_4_9,
input [31:0] ch0_coeff_4_10,
input [31:0] ch1_coeff_1_0,
input [31:0] ch1_coeff_1_1,
input [31:0] ch1_coeff_1_2,
input [31:0] ch1_coeff_1_3,
input [31:0] ch1_coeff_1_4,
input [31:0] ch1_coeff_1_5,
input [31:0] ch1_coeff_1_6,
input [31:0] ch1_coeff_1_7,
input [31:0] ch1_coeff_1_8,
input [31:0] ch1_coeff_1_9,
input [31:0] ch1_coeff_1_10,
input [31:0] ch1_coeff_2_0,
input [31:0] ch1_coeff_2_1,
input [31:0] ch1_coeff_2_2,
input [31:0] ch1_coeff_2_3,
input [31:0] ch1_coeff_2_4,
input [31:0] ch1_coeff_2_5,
input [31:0] ch1_coeff_2_6,
input [31:0] ch1_coeff_2_7,
input [31:0] ch1_coeff_2_8,
input [31:0] ch1_coeff_2_9,
input [31:0] ch1_coeff_2_10,
input [31:0] ch1_coeff_3_0,
input [31:0] ch1_coeff_3_1,
input [31:0] ch1_coeff_3_2,
input [31:0] ch1_coeff_3_3,
input [31:0] ch1_coeff_3_4,
input [31:0] ch1_coeff_3_5,
input [31:0] ch1_coeff_3_6,
input [31:0] ch1_coeff_3_7,
input [31:0] ch1_coeff_3_8,
input [31:0] ch1_coeff_3_9,
input [31:0] ch1_coeff_3_10,
input [31:0] ch1_coeff_4_0,
input [31:0] ch1_coeff_4_1,
input [31:0] ch1_coeff_4_2,
input [31:0] ch1_coeff_4_3,
input [31:0] ch1_coeff_4_4,
input [31:0] ch1_coeff_4_5,
input [31:0] ch1_coeff_4_6,
input [31:0] ch1_coeff_4_7,
input [31:0] ch1_coeff_4_8,
input [31:0] ch1_coeff_4_9,
input [31:0] ch1_coeff_4_10,
input [31:0] ch2_coeff_1_0,
input [31:0] ch2_coeff_1_1,
input [31:0] ch2_coeff_1_2,
input [31:0] ch2_coeff_1_3,
input [31:0] ch2_coeff_1_4,
input [31:0] ch2_coeff_1_5,
input [31:0] ch2_coeff_1_6,
input [31:0] ch2_coeff_1_7,
input [31:0] ch2_coeff_1_8,
input [31:0] ch2_coeff_1_9,
input [31:0] ch2_coeff_1_10,
input [31:0] ch2_coeff_2_0,
input [31:0] ch2_coeff_2_1,
input [31:0] ch2_coeff_2_2,
input [31:0] ch2_coeff_2_3,
input [31:0] ch2_coeff_2_4,
input [31:0] ch2_coeff_2_5,
input [31:0] ch2_coeff_2_6,
input [31:0] ch2_coeff_2_7,
input [31:0] ch2_coeff_2_8,
input [31:0] ch2_coeff_2_9,
input [31:0] ch2_coeff_2_10,
input [31:0] ch2_coeff_3_0,
input [31:0] ch2_coeff_3_1,
input [31:0] ch2_coeff_3_2,
input [31:0] ch2_coeff_3_3,
input [31:0] ch2_coeff_3_4,
input [31:0] ch2_coeff_3_5,
input [31:0] ch2_coeff_3_6,
input [31:0] ch2_coeff_3_7,
input [31:0] ch2_coeff_3_8,
input [31:0] ch2_coeff_3_9,
input [31:0] ch2_coeff_3_10,
input [31:0] ch2_coeff_4_0,
input [31:0] ch2_coeff_4_1,
input [31:0] ch2_coeff_4_2,
input [31:0] ch2_coeff_4_3,
input [31:0] ch2_coeff_4_4,
input [31:0] ch2_coeff_4_5,
input [31:0] ch2_coeff_4_6,
input [31:0] ch2_coeff_4_7,
input [31:0] ch2_coeff_4_8,
input [31:0] ch2_coeff_4_9,
input [31:0] ch2_coeff_4_10,
input [31:0] ch3_coeff_1_0,
input [31:0] ch3_coeff_1_1,
input [31:0] ch3_coeff_1_2,
input [31:0] ch3_coeff_1_3,
input [31:0] ch3_coeff_1_4,
input [31:0] ch3_coeff_1_5,
input [31:0] ch3_coeff_1_6,
input [31:0] ch3_coeff_1_7,
input [31:0] ch3_coeff_1_8,
input [31:0] ch3_coeff_1_9,
input [31:0] ch3_coeff_1_10,
input [31:0] ch3_coeff_2_0,
input [31:0] ch3_coeff_2_1,
input [31:0] ch3_coeff_2_2,
input [31:0] ch3_coeff_2_3,
input [31:0] ch3_coeff_2_4,
input [31:0] ch3_coeff_2_5,
input [31:0] ch3_coeff_2_6,
input [31:0] ch3_coeff_2_7,
input [31:0] ch3_coeff_2_8,
input [31:0] ch3_coeff_2_9,
input [31:0] ch3_coeff_2_10,
input [31:0] ch3_coeff_3_0,
input [31:0] ch3_coeff_3_1,
input [31:0] ch3_coeff_3_2,
input [31:0] ch3_coeff_3_3,
input [31:0] ch3_coeff_3_4,
input [31:0] ch3_coeff_3_5,
input [31:0] ch3_coeff_3_6,
input [31:0] ch3_coeff_3_7,
input [31:0] ch3_coeff_3_8,
input [31:0] ch3_coeff_3_9,
input [31:0] ch3_coeff_3_10,
input [31:0] ch3_coeff_4_0,
input [31:0] ch3_coeff_4_1,
input [31:0] ch3_coeff_4_2,
input [31:0] ch3_coeff_4_3,
input [31:0] ch3_coeff_4_4,
input [31:0] ch3_coeff_4_5,
input [31:0] ch3_coeff_4_6,
input [31:0] ch3_coeff_4_7,
input [31:0] ch3_coeff_4_8,
input [31:0] ch3_coeff_4_9,
input [31:0] ch3_coeff_4_10,
input [31:0] ch4_coeff_1_0,
input [31:0] ch4_coeff_1_1,
input [31:0] ch4_coeff_1_2,
input [31:0] ch4_coeff_1_3,
input [31:0] ch4_coeff_1_4,
input [31:0] ch4_coeff_1_5,
input [31:0] ch4_coeff_1_6,
input [31:0] ch4_coeff_1_7,
input [31:0] ch4_coeff_1_8,
input [31:0] ch4_coeff_1_9,
input [31:0] ch4_coeff_1_10,
input [31:0] ch4_coeff_2_0,
input [31:0] ch4_coeff_2_1,
input [31:0] ch4_coeff_2_2,
input [31:0] ch4_coeff_2_3,
input [31:0] ch4_coeff_2_4,
input [31:0] ch4_coeff_2_5,
input [31:0] ch4_coeff_2_6,
input [31:0] ch4_coeff_2_7,
input [31:0] ch4_coeff_2_8,
input [31:0] ch4_coeff_2_9,
input [31:0] ch4_coeff_2_10,
input [31:0] ch4_coeff_3_0,
input [31:0] ch4_coeff_3_1,
input [31:0] ch4_coeff_3_2,
input [31:0] ch4_coeff_3_3,
input [31:0] ch4_coeff_3_4,
input [31:0] ch4_coeff_3_5,
input [31:0] ch4_coeff_3_6,
input [31:0] ch4_coeff_3_7,
input [31:0] ch4_coeff_3_8,
input [31:0] ch4_coeff_3_9,
input [31:0] ch4_coeff_3_10,
input [31:0] ch4_coeff_4_0,
input [31:0] ch4_coeff_4_1,
input [31:0] ch4_coeff_4_2,
input [31:0] ch4_coeff_4_3,
input [31:0] ch4_coeff_4_4,
input [31:0] ch4_coeff_4_5,
input [31:0] ch4_coeff_4_6,
input [31:0] ch4_coeff_4_7,
input [31:0] ch4_coeff_4_8,
input [31:0] ch4_coeff_4_9,
input [31:0] ch4_coeff_4_10,
input [31:0] ch5_coeff_1_0,
input [31:0] ch5_coeff_1_1,
input [31:0] ch5_coeff_1_2,
input [31:0] ch5_coeff_1_3,
input [31:0] ch5_coeff_1_4,
input [31:0] ch5_coeff_1_5,
input [31:0] ch5_coeff_1_6,
input [31:0] ch5_coeff_1_7,
input [31:0] ch5_coeff_1_8,
input [31:0] ch5_coeff_1_9,
input [31:0] ch5_coeff_1_10,
input [31:0] ch5_coeff_2_0,
input [31:0] ch5_coeff_2_1,
input [31:0] ch5_coeff_2_2,
input [31:0] ch5_coeff_2_3,
input [31:0] ch5_coeff_2_4,
input [31:0] ch5_coeff_2_5,
input [31:0] ch5_coeff_2_6,
input [31:0] ch5_coeff_2_7,
input [31:0] ch5_coeff_2_8,
input [31:0] ch5_coeff_2_9,
input [31:0] ch5_coeff_2_10,
input [31:0] ch5_coeff_3_0,
input [31:0] ch5_coeff_3_1,
input [31:0] ch5_coeff_3_2,
input [31:0] ch5_coeff_3_3,
input [31:0] ch5_coeff_3_4,
input [31:0] ch5_coeff_3_5,
input [31:0] ch5_coeff_3_6,
input [31:0] ch5_coeff_3_7,
input [31:0] ch5_coeff_3_8,
input [31:0] ch5_coeff_3_9,
input [31:0] ch5_coeff_3_10,
input [31:0] ch5_coeff_4_0,
input [31:0] ch5_coeff_4_1,
input [31:0] ch5_coeff_4_2,
input [31:0] ch5_coeff_4_3,
input [31:0] ch5_coeff_4_4,
input [31:0] ch5_coeff_4_5,
input [31:0] ch5_coeff_4_6,
input [31:0] ch5_coeff_4_7,
input [31:0] ch5_coeff_4_8,
input [31:0] ch5_coeff_4_9,
input [31:0] ch5_coeff_4_10,
input [31:0] ch6_coeff_1_0,
input [31:0] ch6_coeff_1_1,
input [31:0] ch6_coeff_1_2,
input [31:0] ch6_coeff_1_3,
input [31:0] ch6_coeff_1_4,
input [31:0] ch6_coeff_1_5,
input [31:0] ch6_coeff_1_6,
input [31:0] ch6_coeff_1_7,
input [31:0] ch6_coeff_1_8,
input [31:0] ch6_coeff_1_9,
input [31:0] ch6_coeff_1_10,
input [31:0] ch6_coeff_2_0,
input [31:0] ch6_coeff_2_1,
input [31:0] ch6_coeff_2_2,
input [31:0] ch6_coeff_2_3,
input [31:0] ch6_coeff_2_4,
input [31:0] ch6_coeff_2_5,
input [31:0] ch6_coeff_2_6,
input [31:0] ch6_coeff_2_7,
input [31:0] ch6_coeff_2_8,
input [31:0] ch6_coeff_2_9,
input [31:0] ch6_coeff_2_10,
input [31:0] ch6_coeff_3_0,
input [31:0] ch6_coeff_3_1,
input [31:0] ch6_coeff_3_2,
input [31:0] ch6_coeff_3_3,
input [31:0] ch6_coeff_3_4,
input [31:0] ch6_coeff_3_5,
input [31:0] ch6_coeff_3_6,
input [31:0] ch6_coeff_3_7,
input [31:0] ch6_coeff_3_8,
input [31:0] ch6_coeff_3_9,
input [31:0] ch6_coeff_3_10,
input [31:0] ch6_coeff_4_0,
input [31:0] ch6_coeff_4_1,
input [31:0] ch6_coeff_4_2,
input [31:0] ch6_coeff_4_3,
input [31:0] ch6_coeff_4_4,
input [31:0] ch6_coeff_4_5,
input [31:0] ch6_coeff_4_6,
input [31:0] ch6_coeff_4_7,
input [31:0] ch6_coeff_4_8,
input [31:0] ch6_coeff_4_9,
input [31:0] ch6_coeff_4_10,
input [31:0] ch7_coeff_1_0,
input [31:0] ch7_coeff_1_1,
input [31:0] ch7_coeff_1_2,
input [31:0] ch7_coeff_1_3,
input [31:0] ch7_coeff_1_4,
input [31:0] ch7_coeff_1_5,
input [31:0] ch7_coeff_1_6,
input [31:0] ch7_coeff_1_7,
input [31:0] ch7_coeff_1_8,
input [31:0] ch7_coeff_1_9,
input [31:0] ch7_coeff_1_10,
input [31:0] ch7_coeff_2_0,
input [31:0] ch7_coeff_2_1,
input [31:0] ch7_coeff_2_2,
input [31:0] ch7_coeff_2_3,
input [31:0] ch7_coeff_2_4,
input [31:0] ch7_coeff_2_5,
input [31:0] ch7_coeff_2_6,
input [31:0] ch7_coeff_2_7,
input [31:0] ch7_coeff_2_8,
input [31:0] ch7_coeff_2_9,
input [31:0] ch7_coeff_2_10,
input [31:0] ch7_coeff_3_0,
input [31:0] ch7_coeff_3_1,
input [31:0] ch7_coeff_3_2,
input [31:0] ch7_coeff_3_3,
input [31:0] ch7_coeff_3_4,
input [31:0] ch7_coeff_3_5,
input [31:0] ch7_coeff_3_6,
input [31:0] ch7_coeff_3_7,
input [31:0] ch7_coeff_3_8,
input [31:0] ch7_coeff_3_9,
input [31:0] ch7_coeff_3_10,
input [31:0] ch7_coeff_4_0,
input [31:0] ch7_coeff_4_1,
input [31:0] ch7_coeff_4_2,
input [31:0] ch7_coeff_4_3,
input [31:0] ch7_coeff_4_4,
input [31:0] ch7_coeff_4_5,
input [31:0] ch7_coeff_4_6,
input [31:0] ch7_coeff_4_7,
input [31:0] ch7_coeff_4_8,
input [31:0] ch7_coeff_4_9,
input [31:0] ch7_coeff_4_10,
input [31:0] ch8_coeff_1_0,
input [31:0] ch8_coeff_1_1,
input [31:0] ch8_coeff_1_2,
input [31:0] ch8_coeff_1_3,
input [31:0] ch8_coeff_1_4,
input [31:0] ch8_coeff_1_5,
input [31:0] ch8_coeff_1_6,
input [31:0] ch8_coeff_1_7,
input [31:0] ch8_coeff_1_8,
input [31:0] ch8_coeff_1_9,
input [31:0] ch8_coeff_1_10,
input [31:0] ch8_coeff_2_0,
input [31:0] ch8_coeff_2_1,
input [31:0] ch8_coeff_2_2,
input [31:0] ch8_coeff_2_3,
input [31:0] ch8_coeff_2_4,
input [31:0] ch8_coeff_2_5,
input [31:0] ch8_coeff_2_6,
input [31:0] ch8_coeff_2_7,
input [31:0] ch8_coeff_2_8,
input [31:0] ch8_coeff_2_9,
input [31:0] ch8_coeff_2_10,
input [31:0] ch8_coeff_3_0,
input [31:0] ch8_coeff_3_1,
input [31:0] ch8_coeff_3_2,
input [31:0] ch8_coeff_3_3,
input [31:0] ch8_coeff_3_4,
input [31:0] ch8_coeff_3_5,
input [31:0] ch8_coeff_3_6,
input [31:0] ch8_coeff_3_7,
input [31:0] ch8_coeff_3_8,
input [31:0] ch8_coeff_3_9,
input [31:0] ch8_coeff_3_10,
input [31:0] ch8_coeff_4_0,
input [31:0] ch8_coeff_4_1,
input [31:0] ch8_coeff_4_2,
input [31:0] ch8_coeff_4_3,
input [31:0] ch8_coeff_4_4,
input [31:0] ch8_coeff_4_5,
input [31:0] ch8_coeff_4_6,
input [31:0] ch8_coeff_4_7,
input [31:0] ch8_coeff_4_8,
input [31:0] ch8_coeff_4_9,
input [31:0] ch8_coeff_4_10,
input [31:0] ch9_coeff_1_0,
input [31:0] ch9_coeff_1_1,
input [31:0] ch9_coeff_1_2,
input [31:0] ch9_coeff_1_3,
input [31:0] ch9_coeff_1_4,
input [31:0] ch9_coeff_1_5,
input [31:0] ch9_coeff_1_6,
input [31:0] ch9_coeff_1_7,
input [31:0] ch9_coeff_1_8,
input [31:0] ch9_coeff_1_9,
input [31:0] ch9_coeff_1_10,
input [31:0] ch9_coeff_2_0,
input [31:0] ch9_coeff_2_1,
input [31:0] ch9_coeff_2_2,
input [31:0] ch9_coeff_2_3,
input [31:0] ch9_coeff_2_4,
input [31:0] ch9_coeff_2_5,
input [31:0] ch9_coeff_2_6,
input [31:0] ch9_coeff_2_7,
input [31:0] ch9_coeff_2_8,
input [31:0] ch9_coeff_2_9,
input [31:0] ch9_coeff_2_10,
input [31:0] ch9_coeff_3_0,
input [31:0] ch9_coeff_3_1,
input [31:0] ch9_coeff_3_2,
input [31:0] ch9_coeff_3_3,
input [31:0] ch9_coeff_3_4,
input [31:0] ch9_coeff_3_5,
input [31:0] ch9_coeff_3_6,
input [31:0] ch9_coeff_3_7,
input [31:0] ch9_coeff_3_8,
input [31:0] ch9_coeff_3_9,
input [31:0] ch9_coeff_3_10,
input [31:0] ch9_coeff_4_0,
input [31:0] ch9_coeff_4_1,
input [31:0] ch9_coeff_4_2,
input [31:0] ch9_coeff_4_3,
input [31:0] ch9_coeff_4_4,
input [31:0] ch9_coeff_4_5,
input [31:0] ch9_coeff_4_6,
input [31:0] ch9_coeff_4_7,
input [31:0] ch9_coeff_4_8,
input [31:0] ch9_coeff_4_9,
input [31:0] ch9_coeff_4_10,
input [31:0] ch10_coeff_1_0,
input [31:0] ch10_coeff_1_1,
input [31:0] ch10_coeff_1_2,
input [31:0] ch10_coeff_1_3,
input [31:0] ch10_coeff_1_4,
input [31:0] ch10_coeff_1_5,
input [31:0] ch10_coeff_1_6,
input [31:0] ch10_coeff_1_7,
input [31:0] ch10_coeff_1_8,
input [31:0] ch10_coeff_1_9,
input [31:0] ch10_coeff_1_10,
input [31:0] ch10_coeff_2_0,
input [31:0] ch10_coeff_2_1,
input [31:0] ch10_coeff_2_2,
input [31:0] ch10_coeff_2_3,
input [31:0] ch10_coeff_2_4,
input [31:0] ch10_coeff_2_5,
input [31:0] ch10_coeff_2_6,
input [31:0] ch10_coeff_2_7,
input [31:0] ch10_coeff_2_8,
input [31:0] ch10_coeff_2_9,
input [31:0] ch10_coeff_2_10,
input [31:0] ch10_coeff_3_0,
input [31:0] ch10_coeff_3_1,
input [31:0] ch10_coeff_3_2,
input [31:0] ch10_coeff_3_3,
input [31:0] ch10_coeff_3_4,
input [31:0] ch10_coeff_3_5,
input [31:0] ch10_coeff_3_6,
input [31:0] ch10_coeff_3_7,
input [31:0] ch10_coeff_3_8,
input [31:0] ch10_coeff_3_9,
input [31:0] ch10_coeff_3_10,
input [31:0] ch10_coeff_4_0,
input [31:0] ch10_coeff_4_1,
input [31:0] ch10_coeff_4_2,
input [31:0] ch10_coeff_4_3,
input [31:0] ch10_coeff_4_4,
input [31:0] ch10_coeff_4_5,
input [31:0] ch10_coeff_4_6,
input [31:0] ch10_coeff_4_7,
input [31:0] ch10_coeff_4_8,
input [31:0] ch10_coeff_4_9,
input [31:0] ch10_coeff_4_10,
input [31:0] ch11_coeff_1_0,
input [31:0] ch11_coeff_1_1,
input [31:0] ch11_coeff_1_2,
input [31:0] ch11_coeff_1_3,
input [31:0] ch11_coeff_1_4,
input [31:0] ch11_coeff_1_5,
input [31:0] ch11_coeff_1_6,
input [31:0] ch11_coeff_1_7,
input [31:0] ch11_coeff_1_8,
input [31:0] ch11_coeff_1_9,
input [31:0] ch11_coeff_1_10,
input [31:0] ch11_coeff_2_0,
input [31:0] ch11_coeff_2_1,
input [31:0] ch11_coeff_2_2,
input [31:0] ch11_coeff_2_3,
input [31:0] ch11_coeff_2_4,
input [31:0] ch11_coeff_2_5,
input [31:0] ch11_coeff_2_6,
input [31:0] ch11_coeff_2_7,
input [31:0] ch11_coeff_2_8,
input [31:0] ch11_coeff_2_9,
input [31:0] ch11_coeff_2_10,
input [31:0] ch11_coeff_3_0,
input [31:0] ch11_coeff_3_1,
input [31:0] ch11_coeff_3_2,
input [31:0] ch11_coeff_3_3,
input [31:0] ch11_coeff_3_4,
input [31:0] ch11_coeff_3_5,
input [31:0] ch11_coeff_3_6,
input [31:0] ch11_coeff_3_7,
input [31:0] ch11_coeff_3_8,
input [31:0] ch11_coeff_3_9,
input [31:0] ch11_coeff_3_10,
input [31:0] ch11_coeff_4_0,
input [31:0] ch11_coeff_4_1,
input [31:0] ch11_coeff_4_2,
input [31:0] ch11_coeff_4_3,
input [31:0] ch11_coeff_4_4,
input [31:0] ch11_coeff_4_5,
input [31:0] ch11_coeff_4_6,
input [31:0] ch11_coeff_4_7,
input [31:0] ch11_coeff_4_8,
input [31:0] ch11_coeff_4_9,
input [31:0] ch11_coeff_4_10,
input [31:0] ch12_coeff_1_0,
input [31:0] ch12_coeff_1_1,
input [31:0] ch12_coeff_1_2,
input [31:0] ch12_coeff_1_3,
input [31:0] ch12_coeff_1_4,
input [31:0] ch12_coeff_1_5,
input [31:0] ch12_coeff_1_6,
input [31:0] ch12_coeff_1_7,
input [31:0] ch12_coeff_1_8,
input [31:0] ch12_coeff_1_9,
input [31:0] ch12_coeff_1_10,
input [31:0] ch12_coeff_2_0,
input [31:0] ch12_coeff_2_1,
input [31:0] ch12_coeff_2_2,
input [31:0] ch12_coeff_2_3,
input [31:0] ch12_coeff_2_4,
input [31:0] ch12_coeff_2_5,
input [31:0] ch12_coeff_2_6,
input [31:0] ch12_coeff_2_7,
input [31:0] ch12_coeff_2_8,
input [31:0] ch12_coeff_2_9,
input [31:0] ch12_coeff_2_10,
input [31:0] ch12_coeff_3_0,
input [31:0] ch12_coeff_3_1,
input [31:0] ch12_coeff_3_2,
input [31:0] ch12_coeff_3_3,
input [31:0] ch12_coeff_3_4,
input [31:0] ch12_coeff_3_5,
input [31:0] ch12_coeff_3_6,
input [31:0] ch12_coeff_3_7,
input [31:0] ch12_coeff_3_8,
input [31:0] ch12_coeff_3_9,
input [31:0] ch12_coeff_3_10,
input [31:0] ch12_coeff_4_0,
input [31:0] ch12_coeff_4_1,
input [31:0] ch12_coeff_4_2,
input [31:0] ch12_coeff_4_3,
input [31:0] ch12_coeff_4_4,
input [31:0] ch12_coeff_4_5,
input [31:0] ch12_coeff_4_6,
input [31:0] ch12_coeff_4_7,
input [31:0] ch12_coeff_4_8,
input [31:0] ch12_coeff_4_9,
input [31:0] ch12_coeff_4_10,
input [31:0] ch13_coeff_1_0,
input [31:0] ch13_coeff_1_1,
input [31:0] ch13_coeff_1_2,
input [31:0] ch13_coeff_1_3,
input [31:0] ch13_coeff_1_4,
input [31:0] ch13_coeff_1_5,
input [31:0] ch13_coeff_1_6,
input [31:0] ch13_coeff_1_7,
input [31:0] ch13_coeff_1_8,
input [31:0] ch13_coeff_1_9,
input [31:0] ch13_coeff_1_10,
input [31:0] ch13_coeff_2_0,
input [31:0] ch13_coeff_2_1,
input [31:0] ch13_coeff_2_2,
input [31:0] ch13_coeff_2_3,
input [31:0] ch13_coeff_2_4,
input [31:0] ch13_coeff_2_5,
input [31:0] ch13_coeff_2_6,
input [31:0] ch13_coeff_2_7,
input [31:0] ch13_coeff_2_8,
input [31:0] ch13_coeff_2_9,
input [31:0] ch13_coeff_2_10,
input [31:0] ch13_coeff_3_0,
input [31:0] ch13_coeff_3_1,
input [31:0] ch13_coeff_3_2,
input [31:0] ch13_coeff_3_3,
input [31:0] ch13_coeff_3_4,
input [31:0] ch13_coeff_3_5,
input [31:0] ch13_coeff_3_6,
input [31:0] ch13_coeff_3_7,
input [31:0] ch13_coeff_3_8,
input [31:0] ch13_coeff_3_9,
input [31:0] ch13_coeff_3_10,
input [31:0] ch13_coeff_4_0,
input [31:0] ch13_coeff_4_1,
input [31:0] ch13_coeff_4_2,
input [31:0] ch13_coeff_4_3,
input [31:0] ch13_coeff_4_4,
input [31:0] ch13_coeff_4_5,
input [31:0] ch13_coeff_4_6,
input [31:0] ch13_coeff_4_7,
input [31:0] ch13_coeff_4_8,
input [31:0] ch13_coeff_4_9,
input [31:0] ch13_coeff_4_10,
input [31:0] ch14_coeff_1_0,
input [31:0] ch14_coeff_1_1,
input [31:0] ch14_coeff_1_2,
input [31:0] ch14_coeff_1_3,
input [31:0] ch14_coeff_1_4,
input [31:0] ch14_coeff_1_5,
input [31:0] ch14_coeff_1_6,
input [31:0] ch14_coeff_1_7,
input [31:0] ch14_coeff_1_8,
input [31:0] ch14_coeff_1_9,
input [31:0] ch14_coeff_1_10,
input [31:0] ch14_coeff_2_0,
input [31:0] ch14_coeff_2_1,
input [31:0] ch14_coeff_2_2,
input [31:0] ch14_coeff_2_3,
input [31:0] ch14_coeff_2_4,
input [31:0] ch14_coeff_2_5,
input [31:0] ch14_coeff_2_6,
input [31:0] ch14_coeff_2_7,
input [31:0] ch14_coeff_2_8,
input [31:0] ch14_coeff_2_9,
input [31:0] ch14_coeff_2_10,
input [31:0] ch14_coeff_3_0,
input [31:0] ch14_coeff_3_1,
input [31:0] ch14_coeff_3_2,
input [31:0] ch14_coeff_3_3,
input [31:0] ch14_coeff_3_4,
input [31:0] ch14_coeff_3_5,
input [31:0] ch14_coeff_3_6,
input [31:0] ch14_coeff_3_7,
input [31:0] ch14_coeff_3_8,
input [31:0] ch14_coeff_3_9,
input [31:0] ch14_coeff_3_10,
input [31:0] ch14_coeff_4_0,
input [31:0] ch14_coeff_4_1,
input [31:0] ch14_coeff_4_2,
input [31:0] ch14_coeff_4_3,
input [31:0] ch14_coeff_4_4,
input [31:0] ch14_coeff_4_5,
input [31:0] ch14_coeff_4_6,
input [31:0] ch14_coeff_4_7,
input [31:0] ch14_coeff_4_8,
input [31:0] ch14_coeff_4_9,
input [31:0] ch14_coeff_4_10,
input [31:0] ch15_coeff_1_0,
input [31:0] ch15_coeff_1_1,
input [31:0] ch15_coeff_1_2,
input [31:0] ch15_coeff_1_3,
input [31:0] ch15_coeff_1_4,
input [31:0] ch15_coeff_1_5,
input [31:0] ch15_coeff_1_6,
input [31:0] ch15_coeff_1_7,
input [31:0] ch15_coeff_1_8,
input [31:0] ch15_coeff_1_9,
input [31:0] ch15_coeff_1_10,
input [31:0] ch15_coeff_2_0,
input [31:0] ch15_coeff_2_1,
input [31:0] ch15_coeff_2_2,
input [31:0] ch15_coeff_2_3,
input [31:0] ch15_coeff_2_4,
input [31:0] ch15_coeff_2_5,
input [31:0] ch15_coeff_2_6,
input [31:0] ch15_coeff_2_7,
input [31:0] ch15_coeff_2_8,
input [31:0] ch15_coeff_2_9,
input [31:0] ch15_coeff_2_10,
input [31:0] ch15_coeff_3_0,
input [31:0] ch15_coeff_3_1,
input [31:0] ch15_coeff_3_2,
input [31:0] ch15_coeff_3_3,
input [31:0] ch15_coeff_3_4,
input [31:0] ch15_coeff_3_5,
input [31:0] ch15_coeff_3_6,
input [31:0] ch15_coeff_3_7,
input [31:0] ch15_coeff_3_8,
input [31:0] ch15_coeff_3_9,
input [31:0] ch15_coeff_3_10,
input [31:0] ch15_coeff_4_0,
input [31:0] ch15_coeff_4_1,
input [31:0] ch15_coeff_4_2,
input [31:0] ch15_coeff_4_3,
input [31:0] ch15_coeff_4_4,
input [31:0] ch15_coeff_4_5,
input [31:0] ch15_coeff_4_6,
input [31:0] ch15_coeff_4_7,
input [31:0] ch15_coeff_4_8,
input [31:0] ch15_coeff_4_9,
input [31:0] ch15_coeff_4_10,
input [31:0] ch16_coeff_1_0,
input [31:0] ch16_coeff_1_1,
input [31:0] ch16_coeff_1_2,
input [31:0] ch16_coeff_1_3,
input [31:0] ch16_coeff_1_4,
input [31:0] ch16_coeff_1_5,
input [31:0] ch16_coeff_1_6,
input [31:0] ch16_coeff_1_7,
input [31:0] ch16_coeff_1_8,
input [31:0] ch16_coeff_1_9,
input [31:0] ch16_coeff_1_10,
input [31:0] ch16_coeff_2_0,
input [31:0] ch16_coeff_2_1,
input [31:0] ch16_coeff_2_2,
input [31:0] ch16_coeff_2_3,
input [31:0] ch16_coeff_2_4,
input [31:0] ch16_coeff_2_5,
input [31:0] ch16_coeff_2_6,
input [31:0] ch16_coeff_2_7,
input [31:0] ch16_coeff_2_8,
input [31:0] ch16_coeff_2_9,
input [31:0] ch16_coeff_2_10,
input [31:0] ch16_coeff_3_0,
input [31:0] ch16_coeff_3_1,
input [31:0] ch16_coeff_3_2,
input [31:0] ch16_coeff_3_3,
input [31:0] ch16_coeff_3_4,
input [31:0] ch16_coeff_3_5,
input [31:0] ch16_coeff_3_6,
input [31:0] ch16_coeff_3_7,
input [31:0] ch16_coeff_3_8,
input [31:0] ch16_coeff_3_9,
input [31:0] ch16_coeff_3_10,
input [31:0] ch16_coeff_4_0,
input [31:0] ch16_coeff_4_1,
input [31:0] ch16_coeff_4_2,
input [31:0] ch16_coeff_4_3,
input [31:0] ch16_coeff_4_4,
input [31:0] ch16_coeff_4_5,
input [31:0] ch16_coeff_4_6,
input [31:0] ch16_coeff_4_7,
input [31:0] ch16_coeff_4_8,
input [31:0] ch16_coeff_4_9,
input [31:0] ch16_coeff_4_10,
input [31:0] ch17_coeff_1_0,
input [31:0] ch17_coeff_1_1,
input [31:0] ch17_coeff_1_2,
input [31:0] ch17_coeff_1_3,
input [31:0] ch17_coeff_1_4,
input [31:0] ch17_coeff_1_5,
input [31:0] ch17_coeff_1_6,
input [31:0] ch17_coeff_1_7,
input [31:0] ch17_coeff_1_8,
input [31:0] ch17_coeff_1_9,
input [31:0] ch17_coeff_1_10,
input [31:0] ch17_coeff_2_0,
input [31:0] ch17_coeff_2_1,
input [31:0] ch17_coeff_2_2,
input [31:0] ch17_coeff_2_3,
input [31:0] ch17_coeff_2_4,
input [31:0] ch17_coeff_2_5,
input [31:0] ch17_coeff_2_6,
input [31:0] ch17_coeff_2_7,
input [31:0] ch17_coeff_2_8,
input [31:0] ch17_coeff_2_9,
input [31:0] ch17_coeff_2_10,
input [31:0] ch17_coeff_3_0,
input [31:0] ch17_coeff_3_1,
input [31:0] ch17_coeff_3_2,
input [31:0] ch17_coeff_3_3,
input [31:0] ch17_coeff_3_4,
input [31:0] ch17_coeff_3_5,
input [31:0] ch17_coeff_3_6,
input [31:0] ch17_coeff_3_7,
input [31:0] ch17_coeff_3_8,
input [31:0] ch17_coeff_3_9,
input [31:0] ch17_coeff_3_10,
input [31:0] ch17_coeff_4_0,
input [31:0] ch17_coeff_4_1,
input [31:0] ch17_coeff_4_2,
input [31:0] ch17_coeff_4_3,
input [31:0] ch17_coeff_4_4,
input [31:0] ch17_coeff_4_5,
input [31:0] ch17_coeff_4_6,
input [31:0] ch17_coeff_4_7,
input [31:0] ch17_coeff_4_8,
input [31:0] ch17_coeff_4_9,
input [31:0] ch17_coeff_4_10,
input [31:0] ch18_coeff_1_0,
input [31:0] ch18_coeff_1_1,
input [31:0] ch18_coeff_1_2,
input [31:0] ch18_coeff_1_3,
input [31:0] ch18_coeff_1_4,
input [31:0] ch18_coeff_1_5,
input [31:0] ch18_coeff_1_6,
input [31:0] ch18_coeff_1_7,
input [31:0] ch18_coeff_1_8,
input [31:0] ch18_coeff_1_9,
input [31:0] ch18_coeff_1_10,
input [31:0] ch18_coeff_2_0,
input [31:0] ch18_coeff_2_1,
input [31:0] ch18_coeff_2_2,
input [31:0] ch18_coeff_2_3,
input [31:0] ch18_coeff_2_4,
input [31:0] ch18_coeff_2_5,
input [31:0] ch18_coeff_2_6,
input [31:0] ch18_coeff_2_7,
input [31:0] ch18_coeff_2_8,
input [31:0] ch18_coeff_2_9,
input [31:0] ch18_coeff_2_10,
input [31:0] ch18_coeff_3_0,
input [31:0] ch18_coeff_3_1,
input [31:0] ch18_coeff_3_2,
input [31:0] ch18_coeff_3_3,
input [31:0] ch18_coeff_3_4,
input [31:0] ch18_coeff_3_5,
input [31:0] ch18_coeff_3_6,
input [31:0] ch18_coeff_3_7,
input [31:0] ch18_coeff_3_8,
input [31:0] ch18_coeff_3_9,
input [31:0] ch18_coeff_3_10,
input [31:0] ch18_coeff_4_0,
input [31:0] ch18_coeff_4_1,
input [31:0] ch18_coeff_4_2,
input [31:0] ch18_coeff_4_3,
input [31:0] ch18_coeff_4_4,
input [31:0] ch18_coeff_4_5,
input [31:0] ch18_coeff_4_6,
input [31:0] ch18_coeff_4_7,
input [31:0] ch18_coeff_4_8,
input [31:0] ch18_coeff_4_9,
input [31:0] ch18_coeff_4_10,
input [31:0] ch19_coeff_1_0,
input [31:0] ch19_coeff_1_1,
input [31:0] ch19_coeff_1_2,
input [31:0] ch19_coeff_1_3,
input [31:0] ch19_coeff_1_4,
input [31:0] ch19_coeff_1_5,
input [31:0] ch19_coeff_1_6,
input [31:0] ch19_coeff_1_7,
input [31:0] ch19_coeff_1_8,
input [31:0] ch19_coeff_1_9,
input [31:0] ch19_coeff_1_10,
input [31:0] ch19_coeff_2_0,
input [31:0] ch19_coeff_2_1,
input [31:0] ch19_coeff_2_2,
input [31:0] ch19_coeff_2_3,
input [31:0] ch19_coeff_2_4,
input [31:0] ch19_coeff_2_5,
input [31:0] ch19_coeff_2_6,
input [31:0] ch19_coeff_2_7,
input [31:0] ch19_coeff_2_8,
input [31:0] ch19_coeff_2_9,
input [31:0] ch19_coeff_2_10,
input [31:0] ch19_coeff_3_0,
input [31:0] ch19_coeff_3_1,
input [31:0] ch19_coeff_3_2,
input [31:0] ch19_coeff_3_3,
input [31:0] ch19_coeff_3_4,
input [31:0] ch19_coeff_3_5,
input [31:0] ch19_coeff_3_6,
input [31:0] ch19_coeff_3_7,
input [31:0] ch19_coeff_3_8,
input [31:0] ch19_coeff_3_9,
input [31:0] ch19_coeff_3_10,
input [31:0] ch19_coeff_4_0,
input [31:0] ch19_coeff_4_1,
input [31:0] ch19_coeff_4_2,
input [31:0] ch19_coeff_4_3,
input [31:0] ch19_coeff_4_4,
input [31:0] ch19_coeff_4_5,
input [31:0] ch19_coeff_4_6,
input [31:0] ch19_coeff_4_7,
input [31:0] ch19_coeff_4_8,
input [31:0] ch19_coeff_4_9,
input [31:0] ch19_coeff_4_10,
input [31:0] ch20_coeff_1_0,
input [31:0] ch20_coeff_1_1,
input [31:0] ch20_coeff_1_2,
input [31:0] ch20_coeff_1_3,
input [31:0] ch20_coeff_1_4,
input [31:0] ch20_coeff_1_5,
input [31:0] ch20_coeff_1_6,
input [31:0] ch20_coeff_1_7,
input [31:0] ch20_coeff_1_8,
input [31:0] ch20_coeff_1_9,
input [31:0] ch20_coeff_1_10,
input [31:0] ch20_coeff_2_0,
input [31:0] ch20_coeff_2_1,
input [31:0] ch20_coeff_2_2,
input [31:0] ch20_coeff_2_3,
input [31:0] ch20_coeff_2_4,
input [31:0] ch20_coeff_2_5,
input [31:0] ch20_coeff_2_6,
input [31:0] ch20_coeff_2_7,
input [31:0] ch20_coeff_2_8,
input [31:0] ch20_coeff_2_9,
input [31:0] ch20_coeff_2_10,
input [31:0] ch20_coeff_3_0,
input [31:0] ch20_coeff_3_1,
input [31:0] ch20_coeff_3_2,
input [31:0] ch20_coeff_3_3,
input [31:0] ch20_coeff_3_4,
input [31:0] ch20_coeff_3_5,
input [31:0] ch20_coeff_3_6,
input [31:0] ch20_coeff_3_7,
input [31:0] ch20_coeff_3_8,
input [31:0] ch20_coeff_3_9,
input [31:0] ch20_coeff_3_10,
input [31:0] ch20_coeff_4_0,
input [31:0] ch20_coeff_4_1,
input [31:0] ch20_coeff_4_2,
input [31:0] ch20_coeff_4_3,
input [31:0] ch20_coeff_4_4,
input [31:0] ch20_coeff_4_5,
input [31:0] ch20_coeff_4_6,
input [31:0] ch20_coeff_4_7,
input [31:0] ch20_coeff_4_8,
input [31:0] ch20_coeff_4_9,
input [31:0] ch20_coeff_4_10,
input [31:0] ch21_coeff_1_0,
input [31:0] ch21_coeff_1_1,
input [31:0] ch21_coeff_1_2,
input [31:0] ch21_coeff_1_3,
input [31:0] ch21_coeff_1_4,
input [31:0] ch21_coeff_1_5,
input [31:0] ch21_coeff_1_6,
input [31:0] ch21_coeff_1_7,
input [31:0] ch21_coeff_1_8,
input [31:0] ch21_coeff_1_9,
input [31:0] ch21_coeff_1_10,
input [31:0] ch21_coeff_2_0,
input [31:0] ch21_coeff_2_1,
input [31:0] ch21_coeff_2_2,
input [31:0] ch21_coeff_2_3,
input [31:0] ch21_coeff_2_4,
input [31:0] ch21_coeff_2_5,
input [31:0] ch21_coeff_2_6,
input [31:0] ch21_coeff_2_7,
input [31:0] ch21_coeff_2_8,
input [31:0] ch21_coeff_2_9,
input [31:0] ch21_coeff_2_10,
input [31:0] ch21_coeff_3_0,
input [31:0] ch21_coeff_3_1,
input [31:0] ch21_coeff_3_2,
input [31:0] ch21_coeff_3_3,
input [31:0] ch21_coeff_3_4,
input [31:0] ch21_coeff_3_5,
input [31:0] ch21_coeff_3_6,
input [31:0] ch21_coeff_3_7,
input [31:0] ch21_coeff_3_8,
input [31:0] ch21_coeff_3_9,
input [31:0] ch21_coeff_3_10,
input [31:0] ch21_coeff_4_0,
input [31:0] ch21_coeff_4_1,
input [31:0] ch21_coeff_4_2,
input [31:0] ch21_coeff_4_3,
input [31:0] ch21_coeff_4_4,
input [31:0] ch21_coeff_4_5,
input [31:0] ch21_coeff_4_6,
input [31:0] ch21_coeff_4_7,
input [31:0] ch21_coeff_4_8,
input [31:0] ch21_coeff_4_9,
input [31:0] ch21_coeff_4_10,
input [31:0] ch22_coeff_1_0,
input [31:0] ch22_coeff_1_1,
input [31:0] ch22_coeff_1_2,
input [31:0] ch22_coeff_1_3,
input [31:0] ch22_coeff_1_4,
input [31:0] ch22_coeff_1_5,
input [31:0] ch22_coeff_1_6,
input [31:0] ch22_coeff_1_7,
input [31:0] ch22_coeff_1_8,
input [31:0] ch22_coeff_1_9,
input [31:0] ch22_coeff_1_10,
input [31:0] ch22_coeff_2_0,
input [31:0] ch22_coeff_2_1,
input [31:0] ch22_coeff_2_2,
input [31:0] ch22_coeff_2_3,
input [31:0] ch22_coeff_2_4,
input [31:0] ch22_coeff_2_5,
input [31:0] ch22_coeff_2_6,
input [31:0] ch22_coeff_2_7,
input [31:0] ch22_coeff_2_8,
input [31:0] ch22_coeff_2_9,
input [31:0] ch22_coeff_2_10,
input [31:0] ch22_coeff_3_0,
input [31:0] ch22_coeff_3_1,
input [31:0] ch22_coeff_3_2,
input [31:0] ch22_coeff_3_3,
input [31:0] ch22_coeff_3_4,
input [31:0] ch22_coeff_3_5,
input [31:0] ch22_coeff_3_6,
input [31:0] ch22_coeff_3_7,
input [31:0] ch22_coeff_3_8,
input [31:0] ch22_coeff_3_9,
input [31:0] ch22_coeff_3_10,
input [31:0] ch22_coeff_4_0,
input [31:0] ch22_coeff_4_1,
input [31:0] ch22_coeff_4_2,
input [31:0] ch22_coeff_4_3,
input [31:0] ch22_coeff_4_4,
input [31:0] ch22_coeff_4_5,
input [31:0] ch22_coeff_4_6,
input [31:0] ch22_coeff_4_7,
input [31:0] ch22_coeff_4_8,
input [31:0] ch22_coeff_4_9,
input [31:0] ch22_coeff_4_10,
input [31:0] ch23_coeff_1_0,
input [31:0] ch23_coeff_1_1,
input [31:0] ch23_coeff_1_2,
input [31:0] ch23_coeff_1_3,
input [31:0] ch23_coeff_1_4,
input [31:0] ch23_coeff_1_5,
input [31:0] ch23_coeff_1_6,
input [31:0] ch23_coeff_1_7,
input [31:0] ch23_coeff_1_8,
input [31:0] ch23_coeff_1_9,
input [31:0] ch23_coeff_1_10,
input [31:0] ch23_coeff_2_0,
input [31:0] ch23_coeff_2_1,
input [31:0] ch23_coeff_2_2,
input [31:0] ch23_coeff_2_3,
input [31:0] ch23_coeff_2_4,
input [31:0] ch23_coeff_2_5,
input [31:0] ch23_coeff_2_6,
input [31:0] ch23_coeff_2_7,
input [31:0] ch23_coeff_2_8,
input [31:0] ch23_coeff_2_9,
input [31:0] ch23_coeff_2_10,
input [31:0] ch23_coeff_3_0,
input [31:0] ch23_coeff_3_1,
input [31:0] ch23_coeff_3_2,
input [31:0] ch23_coeff_3_3,
input [31:0] ch23_coeff_3_4,
input [31:0] ch23_coeff_3_5,
input [31:0] ch23_coeff_3_6,
input [31:0] ch23_coeff_3_7,
input [31:0] ch23_coeff_3_8,
input [31:0] ch23_coeff_3_9,
input [31:0] ch23_coeff_3_10,
input [31:0] ch23_coeff_4_0,
input [31:0] ch23_coeff_4_1,
input [31:0] ch23_coeff_4_2,
input [31:0] ch23_coeff_4_3,
input [31:0] ch23_coeff_4_4,
input [31:0] ch23_coeff_4_5,
input [31:0] ch23_coeff_4_6,
input [31:0] ch23_coeff_4_7,
input [31:0] ch23_coeff_4_8,
input [31:0] ch23_coeff_4_9,
input [31:0] ch23_coeff_4_10,
input [31:0] ch24_coeff_1_0,
input [31:0] ch24_coeff_1_1,
input [31:0] ch24_coeff_1_2,
input [31:0] ch24_coeff_1_3,
input [31:0] ch24_coeff_1_4,
input [31:0] ch24_coeff_1_5,
input [31:0] ch24_coeff_1_6,
input [31:0] ch24_coeff_1_7,
input [31:0] ch24_coeff_1_8,
input [31:0] ch24_coeff_1_9,
input [31:0] ch24_coeff_1_10,
input [31:0] ch24_coeff_2_0,
input [31:0] ch24_coeff_2_1,
input [31:0] ch24_coeff_2_2,
input [31:0] ch24_coeff_2_3,
input [31:0] ch24_coeff_2_4,
input [31:0] ch24_coeff_2_5,
input [31:0] ch24_coeff_2_6,
input [31:0] ch24_coeff_2_7,
input [31:0] ch24_coeff_2_8,
input [31:0] ch24_coeff_2_9,
input [31:0] ch24_coeff_2_10,
input [31:0] ch24_coeff_3_0,
input [31:0] ch24_coeff_3_1,
input [31:0] ch24_coeff_3_2,
input [31:0] ch24_coeff_3_3,
input [31:0] ch24_coeff_3_4,
input [31:0] ch24_coeff_3_5,
input [31:0] ch24_coeff_3_6,
input [31:0] ch24_coeff_3_7,
input [31:0] ch24_coeff_3_8,
input [31:0] ch24_coeff_3_9,
input [31:0] ch24_coeff_3_10,
input [31:0] ch24_coeff_4_0,
input [31:0] ch24_coeff_4_1,
input [31:0] ch24_coeff_4_2,
input [31:0] ch24_coeff_4_3,
input [31:0] ch24_coeff_4_4,
input [31:0] ch24_coeff_4_5,
input [31:0] ch24_coeff_4_6,
input [31:0] ch24_coeff_4_7,
input [31:0] ch24_coeff_4_8,
input [31:0] ch24_coeff_4_9,
input [31:0] ch24_coeff_4_10,
input [31:0] ch25_coeff_1_0,
input [31:0] ch25_coeff_1_1,
input [31:0] ch25_coeff_1_2,
input [31:0] ch25_coeff_1_3,
input [31:0] ch25_coeff_1_4,
input [31:0] ch25_coeff_1_5,
input [31:0] ch25_coeff_1_6,
input [31:0] ch25_coeff_1_7,
input [31:0] ch25_coeff_1_8,
input [31:0] ch25_coeff_1_9,
input [31:0] ch25_coeff_1_10,
input [31:0] ch25_coeff_2_0,
input [31:0] ch25_coeff_2_1,
input [31:0] ch25_coeff_2_2,
input [31:0] ch25_coeff_2_3,
input [31:0] ch25_coeff_2_4,
input [31:0] ch25_coeff_2_5,
input [31:0] ch25_coeff_2_6,
input [31:0] ch25_coeff_2_7,
input [31:0] ch25_coeff_2_8,
input [31:0] ch25_coeff_2_9,
input [31:0] ch25_coeff_2_10,
input [31:0] ch25_coeff_3_0,
input [31:0] ch25_coeff_3_1,
input [31:0] ch25_coeff_3_2,
input [31:0] ch25_coeff_3_3,
input [31:0] ch25_coeff_3_4,
input [31:0] ch25_coeff_3_5,
input [31:0] ch25_coeff_3_6,
input [31:0] ch25_coeff_3_7,
input [31:0] ch25_coeff_3_8,
input [31:0] ch25_coeff_3_9,
input [31:0] ch25_coeff_3_10,
input [31:0] ch25_coeff_4_0,
input [31:0] ch25_coeff_4_1,
input [31:0] ch25_coeff_4_2,
input [31:0] ch25_coeff_4_3,
input [31:0] ch25_coeff_4_4,
input [31:0] ch25_coeff_4_5,
input [31:0] ch25_coeff_4_6,
input [31:0] ch25_coeff_4_7,
input [31:0] ch25_coeff_4_8,
input [31:0] ch25_coeff_4_9,
input [31:0] ch25_coeff_4_10,
input [31:0] ch26_coeff_1_0,
input [31:0] ch26_coeff_1_1,
input [31:0] ch26_coeff_1_2,
input [31:0] ch26_coeff_1_3,
input [31:0] ch26_coeff_1_4,
input [31:0] ch26_coeff_1_5,
input [31:0] ch26_coeff_1_6,
input [31:0] ch26_coeff_1_7,
input [31:0] ch26_coeff_1_8,
input [31:0] ch26_coeff_1_9,
input [31:0] ch26_coeff_1_10,
input [31:0] ch26_coeff_2_0,
input [31:0] ch26_coeff_2_1,
input [31:0] ch26_coeff_2_2,
input [31:0] ch26_coeff_2_3,
input [31:0] ch26_coeff_2_4,
input [31:0] ch26_coeff_2_5,
input [31:0] ch26_coeff_2_6,
input [31:0] ch26_coeff_2_7,
input [31:0] ch26_coeff_2_8,
input [31:0] ch26_coeff_2_9,
input [31:0] ch26_coeff_2_10,
input [31:0] ch26_coeff_3_0,
input [31:0] ch26_coeff_3_1,
input [31:0] ch26_coeff_3_2,
input [31:0] ch26_coeff_3_3,
input [31:0] ch26_coeff_3_4,
input [31:0] ch26_coeff_3_5,
input [31:0] ch26_coeff_3_6,
input [31:0] ch26_coeff_3_7,
input [31:0] ch26_coeff_3_8,
input [31:0] ch26_coeff_3_9,
input [31:0] ch26_coeff_3_10,
input [31:0] ch26_coeff_4_0,
input [31:0] ch26_coeff_4_1,
input [31:0] ch26_coeff_4_2,
input [31:0] ch26_coeff_4_3,
input [31:0] ch26_coeff_4_4,
input [31:0] ch26_coeff_4_5,
input [31:0] ch26_coeff_4_6,
input [31:0] ch26_coeff_4_7,
input [31:0] ch26_coeff_4_8,
input [31:0] ch26_coeff_4_9,
input [31:0] ch26_coeff_4_10,
input [31:0] ch27_coeff_1_0,
input [31:0] ch27_coeff_1_1,
input [31:0] ch27_coeff_1_2,
input [31:0] ch27_coeff_1_3,
input [31:0] ch27_coeff_1_4,
input [31:0] ch27_coeff_1_5,
input [31:0] ch27_coeff_1_6,
input [31:0] ch27_coeff_1_7,
input [31:0] ch27_coeff_1_8,
input [31:0] ch27_coeff_1_9,
input [31:0] ch27_coeff_1_10,
input [31:0] ch27_coeff_2_0,
input [31:0] ch27_coeff_2_1,
input [31:0] ch27_coeff_2_2,
input [31:0] ch27_coeff_2_3,
input [31:0] ch27_coeff_2_4,
input [31:0] ch27_coeff_2_5,
input [31:0] ch27_coeff_2_6,
input [31:0] ch27_coeff_2_7,
input [31:0] ch27_coeff_2_8,
input [31:0] ch27_coeff_2_9,
input [31:0] ch27_coeff_2_10,
input [31:0] ch27_coeff_3_0,
input [31:0] ch27_coeff_3_1,
input [31:0] ch27_coeff_3_2,
input [31:0] ch27_coeff_3_3,
input [31:0] ch27_coeff_3_4,
input [31:0] ch27_coeff_3_5,
input [31:0] ch27_coeff_3_6,
input [31:0] ch27_coeff_3_7,
input [31:0] ch27_coeff_3_8,
input [31:0] ch27_coeff_3_9,
input [31:0] ch27_coeff_3_10,
input [31:0] ch27_coeff_4_0,
input [31:0] ch27_coeff_4_1,
input [31:0] ch27_coeff_4_2,
input [31:0] ch27_coeff_4_3,
input [31:0] ch27_coeff_4_4,
input [31:0] ch27_coeff_4_5,
input [31:0] ch27_coeff_4_6,
input [31:0] ch27_coeff_4_7,
input [31:0] ch27_coeff_4_8,
input [31:0] ch27_coeff_4_9,
input [31:0] ch27_coeff_4_10,
input [31:0] ch28_coeff_1_0,
input [31:0] ch28_coeff_1_1,
input [31:0] ch28_coeff_1_2,
input [31:0] ch28_coeff_1_3,
input [31:0] ch28_coeff_1_4,
input [31:0] ch28_coeff_1_5,
input [31:0] ch28_coeff_1_6,
input [31:0] ch28_coeff_1_7,
input [31:0] ch28_coeff_1_8,
input [31:0] ch28_coeff_1_9,
input [31:0] ch28_coeff_1_10,
input [31:0] ch28_coeff_2_0,
input [31:0] ch28_coeff_2_1,
input [31:0] ch28_coeff_2_2,
input [31:0] ch28_coeff_2_3,
input [31:0] ch28_coeff_2_4,
input [31:0] ch28_coeff_2_5,
input [31:0] ch28_coeff_2_6,
input [31:0] ch28_coeff_2_7,
input [31:0] ch28_coeff_2_8,
input [31:0] ch28_coeff_2_9,
input [31:0] ch28_coeff_2_10,
input [31:0] ch28_coeff_3_0,
input [31:0] ch28_coeff_3_1,
input [31:0] ch28_coeff_3_2,
input [31:0] ch28_coeff_3_3,
input [31:0] ch28_coeff_3_4,
input [31:0] ch28_coeff_3_5,
input [31:0] ch28_coeff_3_6,
input [31:0] ch28_coeff_3_7,
input [31:0] ch28_coeff_3_8,
input [31:0] ch28_coeff_3_9,
input [31:0] ch28_coeff_3_10,
input [31:0] ch28_coeff_4_0,
input [31:0] ch28_coeff_4_1,
input [31:0] ch28_coeff_4_2,
input [31:0] ch28_coeff_4_3,
input [31:0] ch28_coeff_4_4,
input [31:0] ch28_coeff_4_5,
input [31:0] ch28_coeff_4_6,
input [31:0] ch28_coeff_4_7,
input [31:0] ch28_coeff_4_8,
input [31:0] ch28_coeff_4_9,
input [31:0] ch28_coeff_4_10,
input [31:0] ch29_coeff_1_0,
input [31:0] ch29_coeff_1_1,
input [31:0] ch29_coeff_1_2,
input [31:0] ch29_coeff_1_3,
input [31:0] ch29_coeff_1_4,
input [31:0] ch29_coeff_1_5,
input [31:0] ch29_coeff_1_6,
input [31:0] ch29_coeff_1_7,
input [31:0] ch29_coeff_1_8,
input [31:0] ch29_coeff_1_9,
input [31:0] ch29_coeff_1_10,
input [31:0] ch29_coeff_2_0,
input [31:0] ch29_coeff_2_1,
input [31:0] ch29_coeff_2_2,
input [31:0] ch29_coeff_2_3,
input [31:0] ch29_coeff_2_4,
input [31:0] ch29_coeff_2_5,
input [31:0] ch29_coeff_2_6,
input [31:0] ch29_coeff_2_7,
input [31:0] ch29_coeff_2_8,
input [31:0] ch29_coeff_2_9,
input [31:0] ch29_coeff_2_10,
input [31:0] ch29_coeff_3_0,
input [31:0] ch29_coeff_3_1,
input [31:0] ch29_coeff_3_2,
input [31:0] ch29_coeff_3_3,
input [31:0] ch29_coeff_3_4,
input [31:0] ch29_coeff_3_5,
input [31:0] ch29_coeff_3_6,
input [31:0] ch29_coeff_3_7,
input [31:0] ch29_coeff_3_8,
input [31:0] ch29_coeff_3_9,
input [31:0] ch29_coeff_3_10,
input [31:0] ch29_coeff_4_0,
input [31:0] ch29_coeff_4_1,
input [31:0] ch29_coeff_4_2,
input [31:0] ch29_coeff_4_3,
input [31:0] ch29_coeff_4_4,
input [31:0] ch29_coeff_4_5,
input [31:0] ch29_coeff_4_6,
input [31:0] ch29_coeff_4_7,
input [31:0] ch29_coeff_4_8,
input [31:0] ch29_coeff_4_9,
input [31:0] ch29_coeff_4_10,
input [31:0] ch30_coeff_1_0,
input [31:0] ch30_coeff_1_1,
input [31:0] ch30_coeff_1_2,
input [31:0] ch30_coeff_1_3,
input [31:0] ch30_coeff_1_4,
input [31:0] ch30_coeff_1_5,
input [31:0] ch30_coeff_1_6,
input [31:0] ch30_coeff_1_7,
input [31:0] ch30_coeff_1_8,
input [31:0] ch30_coeff_1_9,
input [31:0] ch30_coeff_1_10,
input [31:0] ch30_coeff_2_0,
input [31:0] ch30_coeff_2_1,
input [31:0] ch30_coeff_2_2,
input [31:0] ch30_coeff_2_3,
input [31:0] ch30_coeff_2_4,
input [31:0] ch30_coeff_2_5,
input [31:0] ch30_coeff_2_6,
input [31:0] ch30_coeff_2_7,
input [31:0] ch30_coeff_2_8,
input [31:0] ch30_coeff_2_9,
input [31:0] ch30_coeff_2_10,
input [31:0] ch30_coeff_3_0,
input [31:0] ch30_coeff_3_1,
input [31:0] ch30_coeff_3_2,
input [31:0] ch30_coeff_3_3,
input [31:0] ch30_coeff_3_4,
input [31:0] ch30_coeff_3_5,
input [31:0] ch30_coeff_3_6,
input [31:0] ch30_coeff_3_7,
input [31:0] ch30_coeff_3_8,
input [31:0] ch30_coeff_3_9,
input [31:0] ch30_coeff_3_10,
input [31:0] ch30_coeff_4_0,
input [31:0] ch30_coeff_4_1,
input [31:0] ch30_coeff_4_2,
input [31:0] ch30_coeff_4_3,
input [31:0] ch30_coeff_4_4,
input [31:0] ch30_coeff_4_5,
input [31:0] ch30_coeff_4_6,
input [31:0] ch30_coeff_4_7,
input [31:0] ch30_coeff_4_8,
input [31:0] ch30_coeff_4_9,
input [31:0] ch30_coeff_4_10,
input [31:0] ch31_coeff_1_0,
input [31:0] ch31_coeff_1_1,
input [31:0] ch31_coeff_1_2,
input [31:0] ch31_coeff_1_3,
input [31:0] ch31_coeff_1_4,
input [31:0] ch31_coeff_1_5,
input [31:0] ch31_coeff_1_6,
input [31:0] ch31_coeff_1_7,
input [31:0] ch31_coeff_1_8,
input [31:0] ch31_coeff_1_9,
input [31:0] ch31_coeff_1_10,
input [31:0] ch31_coeff_2_0,
input [31:0] ch31_coeff_2_1,
input [31:0] ch31_coeff_2_2,
input [31:0] ch31_coeff_2_3,
input [31:0] ch31_coeff_2_4,
input [31:0] ch31_coeff_2_5,
input [31:0] ch31_coeff_2_6,
input [31:0] ch31_coeff_2_7,
input [31:0] ch31_coeff_2_8,
input [31:0] ch31_coeff_2_9,
input [31:0] ch31_coeff_2_10,
input [31:0] ch31_coeff_3_0,
input [31:0] ch31_coeff_3_1,
input [31:0] ch31_coeff_3_2,
input [31:0] ch31_coeff_3_3,
input [31:0] ch31_coeff_3_4,
input [31:0] ch31_coeff_3_5,
input [31:0] ch31_coeff_3_6,
input [31:0] ch31_coeff_3_7,
input [31:0] ch31_coeff_3_8,
input [31:0] ch31_coeff_3_9,
input [31:0] ch31_coeff_3_10,
input [31:0] ch31_coeff_4_0,
input [31:0] ch31_coeff_4_1,
input [31:0] ch31_coeff_4_2,
input [31:0] ch31_coeff_4_3,
input [31:0] ch31_coeff_4_4,
input [31:0] ch31_coeff_4_5,
input [31:0] ch31_coeff_4_6,
input [31:0] ch31_coeff_4_7,
input [31:0] ch31_coeff_4_8,
input [31:0] ch31_coeff_4_9,
input [31:0] ch31_coeff_4_10,
input [31:0] ch0_neg_mean_1,
input [31:0] ch0_recip_stdev_1,
input [31:0] ch0_neg_mean_2,
input [31:0] ch0_recip_stdev_2,
input [31:0] ch0_neg_mean_3,
input [31:0] ch0_recip_stdev_3,
input [31:0] ch0_neg_mean_4,
input [31:0] ch0_recip_stdev_4,
input [31:0] ch1_neg_mean_1,
input [31:0] ch1_recip_stdev_1,
input [31:0] ch1_neg_mean_2,
input [31:0] ch1_recip_stdev_2,
input [31:0] ch1_neg_mean_3,
input [31:0] ch1_recip_stdev_3,
input [31:0] ch1_neg_mean_4,
input [31:0] ch1_recip_stdev_4,
input [31:0] ch2_neg_mean_1,
input [31:0] ch2_recip_stdev_1,
input [31:0] ch2_neg_mean_2,
input [31:0] ch2_recip_stdev_2,
input [31:0] ch2_neg_mean_3,
input [31:0] ch2_recip_stdev_3,
input [31:0] ch2_neg_mean_4,
input [31:0] ch2_recip_stdev_4,
input [31:0] ch3_neg_mean_1,
input [31:0] ch3_recip_stdev_1,
input [31:0] ch3_neg_mean_2,
input [31:0] ch3_recip_stdev_2,
input [31:0] ch3_neg_mean_3,
input [31:0] ch3_recip_stdev_3,
input [31:0] ch3_neg_mean_4,
input [31:0] ch3_recip_stdev_4,
input [31:0] ch4_neg_mean_1,
input [31:0] ch4_recip_stdev_1,
input [31:0] ch4_neg_mean_2,
input [31:0] ch4_recip_stdev_2,
input [31:0] ch4_neg_mean_3,
input [31:0] ch4_recip_stdev_3,
input [31:0] ch4_neg_mean_4,
input [31:0] ch4_recip_stdev_4,
input [31:0] ch5_neg_mean_1,
input [31:0] ch5_recip_stdev_1,
input [31:0] ch5_neg_mean_2,
input [31:0] ch5_recip_stdev_2,
input [31:0] ch5_neg_mean_3,
input [31:0] ch5_recip_stdev_3,
input [31:0] ch5_neg_mean_4,
input [31:0] ch5_recip_stdev_4,
input [31:0] ch6_neg_mean_1,
input [31:0] ch6_recip_stdev_1,
input [31:0] ch6_neg_mean_2,
input [31:0] ch6_recip_stdev_2,
input [31:0] ch6_neg_mean_3,
input [31:0] ch6_recip_stdev_3,
input [31:0] ch6_neg_mean_4,
input [31:0] ch6_recip_stdev_4,
input [31:0] ch7_neg_mean_1,
input [31:0] ch7_recip_stdev_1,
input [31:0] ch7_neg_mean_2,
input [31:0] ch7_recip_stdev_2,
input [31:0] ch7_neg_mean_3,
input [31:0] ch7_recip_stdev_3,
input [31:0] ch7_neg_mean_4,
input [31:0] ch7_recip_stdev_4,
input [31:0] ch8_neg_mean_1,
input [31:0] ch8_recip_stdev_1,
input [31:0] ch8_neg_mean_2,
input [31:0] ch8_recip_stdev_2,
input [31:0] ch8_neg_mean_3,
input [31:0] ch8_recip_stdev_3,
input [31:0] ch8_neg_mean_4,
input [31:0] ch8_recip_stdev_4,
input [31:0] ch9_neg_mean_1,
input [31:0] ch9_recip_stdev_1,
input [31:0] ch9_neg_mean_2,
input [31:0] ch9_recip_stdev_2,
input [31:0] ch9_neg_mean_3,
input [31:0] ch9_recip_stdev_3,
input [31:0] ch9_neg_mean_4,
input [31:0] ch9_recip_stdev_4,
input [31:0] ch10_neg_mean_1,
input [31:0] ch10_recip_stdev_1,
input [31:0] ch10_neg_mean_2,
input [31:0] ch10_recip_stdev_2,
input [31:0] ch10_neg_mean_3,
input [31:0] ch10_recip_stdev_3,
input [31:0] ch10_neg_mean_4,
input [31:0] ch10_recip_stdev_4,
input [31:0] ch11_neg_mean_1,
input [31:0] ch11_recip_stdev_1,
input [31:0] ch11_neg_mean_2,
input [31:0] ch11_recip_stdev_2,
input [31:0] ch11_neg_mean_3,
input [31:0] ch11_recip_stdev_3,
input [31:0] ch11_neg_mean_4,
input [31:0] ch11_recip_stdev_4,
input [31:0] ch12_neg_mean_1,
input [31:0] ch12_recip_stdev_1,
input [31:0] ch12_neg_mean_2,
input [31:0] ch12_recip_stdev_2,
input [31:0] ch12_neg_mean_3,
input [31:0] ch12_recip_stdev_3,
input [31:0] ch12_neg_mean_4,
input [31:0] ch12_recip_stdev_4,
input [31:0] ch13_neg_mean_1,
input [31:0] ch13_recip_stdev_1,
input [31:0] ch13_neg_mean_2,
input [31:0] ch13_recip_stdev_2,
input [31:0] ch13_neg_mean_3,
input [31:0] ch13_recip_stdev_3,
input [31:0] ch13_neg_mean_4,
input [31:0] ch13_recip_stdev_4,
input [31:0] ch14_neg_mean_1,
input [31:0] ch14_recip_stdev_1,
input [31:0] ch14_neg_mean_2,
input [31:0] ch14_recip_stdev_2,
input [31:0] ch14_neg_mean_3,
input [31:0] ch14_recip_stdev_3,
input [31:0] ch14_neg_mean_4,
input [31:0] ch14_recip_stdev_4,
input [31:0] ch15_neg_mean_1,
input [31:0] ch15_recip_stdev_1,
input [31:0] ch15_neg_mean_2,
input [31:0] ch15_recip_stdev_2,
input [31:0] ch15_neg_mean_3,
input [31:0] ch15_recip_stdev_3,
input [31:0] ch15_neg_mean_4,
input [31:0] ch15_recip_stdev_4,
input [31:0] ch16_neg_mean_1,
input [31:0] ch16_recip_stdev_1,
input [31:0] ch16_neg_mean_2,
input [31:0] ch16_recip_stdev_2,
input [31:0] ch16_neg_mean_3,
input [31:0] ch16_recip_stdev_3,
input [31:0] ch16_neg_mean_4,
input [31:0] ch16_recip_stdev_4,
input [31:0] ch17_neg_mean_1,
input [31:0] ch17_recip_stdev_1,
input [31:0] ch17_neg_mean_2,
input [31:0] ch17_recip_stdev_2,
input [31:0] ch17_neg_mean_3,
input [31:0] ch17_recip_stdev_3,
input [31:0] ch17_neg_mean_4,
input [31:0] ch17_recip_stdev_4,
input [31:0] ch18_neg_mean_1,
input [31:0] ch18_recip_stdev_1,
input [31:0] ch18_neg_mean_2,
input [31:0] ch18_recip_stdev_2,
input [31:0] ch18_neg_mean_3,
input [31:0] ch18_recip_stdev_3,
input [31:0] ch18_neg_mean_4,
input [31:0] ch18_recip_stdev_4,
input [31:0] ch19_neg_mean_1,
input [31:0] ch19_recip_stdev_1,
input [31:0] ch19_neg_mean_2,
input [31:0] ch19_recip_stdev_2,
input [31:0] ch19_neg_mean_3,
input [31:0] ch19_recip_stdev_3,
input [31:0] ch19_neg_mean_4,
input [31:0] ch19_recip_stdev_4,
input [31:0] ch20_neg_mean_1,
input [31:0] ch20_recip_stdev_1,
input [31:0] ch20_neg_mean_2,
input [31:0] ch20_recip_stdev_2,
input [31:0] ch20_neg_mean_3,
input [31:0] ch20_recip_stdev_3,
input [31:0] ch20_neg_mean_4,
input [31:0] ch20_recip_stdev_4,
input [31:0] ch21_neg_mean_1,
input [31:0] ch21_recip_stdev_1,
input [31:0] ch21_neg_mean_2,
input [31:0] ch21_recip_stdev_2,
input [31:0] ch21_neg_mean_3,
input [31:0] ch21_recip_stdev_3,
input [31:0] ch21_neg_mean_4,
input [31:0] ch21_recip_stdev_4,
input [31:0] ch22_neg_mean_1,
input [31:0] ch22_recip_stdev_1,
input [31:0] ch22_neg_mean_2,
input [31:0] ch22_recip_stdev_2,
input [31:0] ch22_neg_mean_3,
input [31:0] ch22_recip_stdev_3,
input [31:0] ch22_neg_mean_4,
input [31:0] ch22_recip_stdev_4,
input [31:0] ch23_neg_mean_1,
input [31:0] ch23_recip_stdev_1,
input [31:0] ch23_neg_mean_2,
input [31:0] ch23_recip_stdev_2,
input [31:0] ch23_neg_mean_3,
input [31:0] ch23_recip_stdev_3,
input [31:0] ch23_neg_mean_4,
input [31:0] ch23_recip_stdev_4,
input [31:0] ch24_neg_mean_1,
input [31:0] ch24_recip_stdev_1,
input [31:0] ch24_neg_mean_2,
input [31:0] ch24_recip_stdev_2,
input [31:0] ch24_neg_mean_3,
input [31:0] ch24_recip_stdev_3,
input [31:0] ch24_neg_mean_4,
input [31:0] ch24_recip_stdev_4,
input [31:0] ch25_neg_mean_1,
input [31:0] ch25_recip_stdev_1,
input [31:0] ch25_neg_mean_2,
input [31:0] ch25_recip_stdev_2,
input [31:0] ch25_neg_mean_3,
input [31:0] ch25_recip_stdev_3,
input [31:0] ch25_neg_mean_4,
input [31:0] ch25_recip_stdev_4,
input [31:0] ch26_neg_mean_1,
input [31:0] ch26_recip_stdev_1,
input [31:0] ch26_neg_mean_2,
input [31:0] ch26_recip_stdev_2,
input [31:0] ch26_neg_mean_3,
input [31:0] ch26_recip_stdev_3,
input [31:0] ch26_neg_mean_4,
input [31:0] ch26_recip_stdev_4,
input [31:0] ch27_neg_mean_1,
input [31:0] ch27_recip_stdev_1,
input [31:0] ch27_neg_mean_2,
input [31:0] ch27_recip_stdev_2,
input [31:0] ch27_neg_mean_3,
input [31:0] ch27_recip_stdev_3,
input [31:0] ch27_neg_mean_4,
input [31:0] ch27_recip_stdev_4,
input [31:0] ch28_neg_mean_1,
input [31:0] ch28_recip_stdev_1,
input [31:0] ch28_neg_mean_2,
input [31:0] ch28_recip_stdev_2,
input [31:0] ch28_neg_mean_3,
input [31:0] ch28_recip_stdev_3,
input [31:0] ch28_neg_mean_4,
input [31:0] ch28_recip_stdev_4,
input [31:0] ch29_neg_mean_1,
input [31:0] ch29_recip_stdev_1,
input [31:0] ch29_neg_mean_2,
input [31:0] ch29_recip_stdev_2,
input [31:0] ch29_neg_mean_3,
input [31:0] ch29_recip_stdev_3,
input [31:0] ch29_neg_mean_4,
input [31:0] ch29_recip_stdev_4,
input [31:0] ch30_neg_mean_1,
input [31:0] ch30_recip_stdev_1,
input [31:0] ch30_neg_mean_2,
input [31:0] ch30_recip_stdev_2,
input [31:0] ch30_neg_mean_3,
input [31:0] ch30_recip_stdev_3,
input [31:0] ch30_neg_mean_4,
input [31:0] ch30_recip_stdev_4,
input [31:0] ch31_neg_mean_1,
input [31:0] ch31_recip_stdev_1,
input [31:0] ch31_neg_mean_2,
input [31:0] ch31_recip_stdev_2,
input [31:0] ch31_neg_mean_3,
input [31:0] ch31_recip_stdev_3,
input [31:0] ch31_neg_mean_4,
input [31:0] ch31_recip_stdev_4,
input clk,
input reset,
output srdyo, 
input srdyi, 
input [20:0] ch0_x_adc,
output [20:0] ch0_x_lin,
input [19:0] ch0_section_limit,
input [20:0] ch1_x_adc,
output [20:0] ch1_x_lin,
input [19:0] ch1_section_limit,
input [20:0] ch2_x_adc,
output [20:0] ch2_x_lin,
input [19:0] ch2_section_limit,
input [20:0] ch3_x_adc,
output [20:0] ch3_x_lin,
input [19:0] ch3_section_limit,
input [20:0] ch4_x_adc,
output [20:0] ch4_x_lin,
input [19:0] ch4_section_limit,
input [20:0] ch5_x_adc,
output [20:0] ch5_x_lin,
input [19:0] ch5_section_limit,
input [20:0] ch6_x_adc,
output [20:0] ch6_x_lin,
input [19:0] ch6_section_limit,
input [20:0] ch7_x_adc,
output [20:0] ch7_x_lin,
input [19:0] ch7_section_limit,
input [20:0] ch8_x_adc,
output [20:0] ch8_x_lin,
input [19:0] ch8_section_limit,
input [20:0] ch9_x_adc,
output [20:0] ch9_x_lin,
input [19:0] ch9_section_limit,
input [20:0] ch10_x_adc,
output [20:0] ch10_x_lin,
input [19:0] ch10_section_limit,
input [20:0] ch11_x_adc,
output [20:0] ch11_x_lin,
input [19:0] ch11_section_limit,
input [20:0] ch12_x_adc,
output [20:0] ch12_x_lin,
input [19:0] ch12_section_limit,
input [20:0] ch13_x_adc,
output [20:0] ch13_x_lin,
input [19:0] ch13_section_limit,
input [20:0] ch14_x_adc,
output [20:0] ch14_x_lin,
input [19:0] ch14_section_limit,
input [20:0] ch15_x_adc,
output [20:0] ch15_x_lin,
input [19:0] ch15_section_limit,
input [20:0] ch16_x_adc,
output [20:0] ch16_x_lin,
input [19:0] ch16_section_limit,
input [20:0] ch17_x_adc,
output [20:0] ch17_x_lin,
input [19:0] ch17_section_limit,
input [20:0] ch18_x_adc,
output [20:0] ch18_x_lin,
input [19:0] ch18_section_limit,
input [20:0] ch19_x_adc,
output [20:0] ch19_x_lin,
input [19:0] ch19_section_limit,
input [20:0] ch20_x_adc,
output [20:0] ch20_x_lin,
input [19:0] ch20_section_limit,
input [20:0] ch21_x_adc,
output [20:0] ch21_x_lin,
input [19:0] ch21_section_limit,
input [20:0] ch22_x_adc,
output [20:0] ch22_x_lin,
input [19:0] ch22_section_limit,
input [20:0] ch23_x_adc,
output [20:0] ch23_x_lin,
input [19:0] ch23_section_limit,
input [20:0] ch24_x_adc,
output [20:0] ch24_x_lin,
input [19:0] ch24_section_limit,
input [20:0] ch25_x_adc,
output [20:0] ch25_x_lin,
input [19:0] ch25_section_limit,
input [20:0] ch26_x_adc,
output [20:0] ch26_x_lin,
input [19:0] ch26_section_limit,
input [20:0] ch27_x_adc,
output [20:0] ch27_x_lin,
input [19:0] ch27_section_limit,
input [20:0] ch28_x_adc,
output [20:0] ch28_x_lin,
input [19:0] ch28_section_limit,
input [20:0] ch29_x_adc,
output [20:0] ch29_x_lin,
input [19:0] ch29_section_limit,
input [20:0] ch30_x_adc,
output [20:0] ch30_x_lin,
input [19:0] ch30_section_limit,
input [20:0] ch31_x_adc,
output [20:0] ch31_x_lin,
input [19:0] ch31_section_limit
);


wire [15:0] section_select;
wire [20:0] buffer_out;
wire srdyi_buffer;
wire srdyo_NLC1ch;
wire [20:0] fp_res;
wire del;

delay d(.clk(clk), .reset(reset), .enable(srdyo_NLC1ch), .del(del));


buffer_inputs b (.clk(clk), .reset(reset), .srdyi_1(srdyi), .srdyi_2(del),
  .fp_input_0(ch0_x_adc), .ch0_section_limit(ch0_section_limit), 
  .fp_input_1(ch1_x_adc), .ch1_section_limit(ch1_section_limit), 
  .fp_input_2(ch2_x_adc), .ch2_section_limit(ch2_section_limit), 
  .fp_input_3(ch3_x_adc), .ch3_section_limit(ch3_section_limit), 
  .fp_input_4(ch4_x_adc), .ch4_section_limit(ch4_section_limit), 
  .fp_input_5(ch5_x_adc), .ch5_section_limit(ch5_section_limit), 
  .fp_input_6(ch6_x_adc), .ch6_section_limit(ch6_section_limit), 
  .fp_input_7(ch7_x_adc), .ch7_section_limit(ch7_section_limit), 
  .fp_input_8(ch8_x_adc), .ch8_section_limit(ch8_section_limit), 
  .fp_input_9(ch9_x_adc), .ch9_section_limit(ch9_section_limit), 
  .fp_input_10(ch10_x_adc), .ch10_section_limit(ch10_section_limit), 
  .fp_input_11(ch11_x_adc), .ch11_section_limit(ch11_section_limit), 
  .fp_input_12(ch12_x_adc), .ch12_section_limit(ch12_section_limit), 
  .fp_input_13(ch13_x_adc), .ch13_section_limit(ch13_section_limit), 
  .fp_input_14(ch14_x_adc), .ch14_section_limit(ch14_section_limit), 
  .fp_input_15(ch15_x_adc), .ch15_section_limit(ch15_section_limit), 
  .fp_input_16(ch16_x_adc), .ch16_section_limit(ch16_section_limit), 
  .fp_input_17(ch17_x_adc), .ch17_section_limit(ch17_section_limit), 
  .fp_input_18(ch18_x_adc), .ch18_section_limit(ch18_section_limit), 
  .fp_input_19(ch19_x_adc), .ch19_section_limit(ch19_section_limit), 
  .fp_input_20(ch20_x_adc), .ch20_section_limit(ch20_section_limit), 
  .fp_input_21(ch21_x_adc), .ch21_section_limit(ch21_section_limit), 
  .fp_input_22(ch22_x_adc), .ch22_section_limit(ch22_section_limit), 
  .fp_input_23(ch23_x_adc), .ch23_section_limit(ch23_section_limit), 
  .fp_input_24(ch24_x_adc), .ch24_section_limit(ch24_section_limit), 
  .fp_input_25(ch25_x_adc), .ch25_section_limit(ch25_section_limit), 
  .fp_input_26(ch26_x_adc), .ch26_section_limit(ch26_section_limit), 
  .fp_input_27(ch27_x_adc), .ch27_section_limit(ch27_section_limit), 
  .fp_input_28(ch28_x_adc), .ch28_section_limit(ch28_section_limit), 
  .fp_input_29(ch29_x_adc), .ch29_section_limit(ch29_section_limit), 
  .fp_input_30(ch30_x_adc), .ch30_section_limit(ch30_section_limit), 
  .fp_input_31(ch31_x_adc), .ch31_section_limit(ch31_section_limit),
  .section_select(section_select), .out(buffer_out), .srdyo(srdyo_buffer));

NLC_1ch NLC (.clk(clk),.reset(reset),.srdyi(srdyo_buffer),.srdyo(srdyo_NLC1ch),.x_adc(buffer_out),
	.x_lin(fp_res),.recip_stdev_1(ch0_recip_stdev_1),
	.recip_stdev_2(ch0_recip_stdev_2),.recip_stdev_3(ch0_recip_stdev_3),.recip_stdev_4(ch0_recip_stdev_4),
	.neg_mean_1(ch0_neg_mean_1),.neg_mean_2(ch0_neg_mean_2),.neg_mean_3(ch0_neg_mean_3),
	.neg_mean_4(ch0_neg_mean_4),
	.coeff_1_0(ch0_coeff_1_0),.coeff_1_1(ch0_coeff_1_1),.coeff_1_2(ch0_coeff_1_2),.coeff_1_3(ch0_coeff_1_3),
	.coeff_1_4(ch0_coeff_1_4),.coeff_1_5(ch0_coeff_1_5),
	.coeff_1_6(ch0_coeff_1_6),.coeff_1_7(ch0_coeff_1_7),.coeff_1_8(ch0_coeff_1_8),.coeff_1_9(ch0_coeff_1_9),
	.coeff_1_10(ch0_coeff_1_10),.coeff_2_0(ch0_coeff_2_0),
	.coeff_2_1(ch0_coeff_2_1),.coeff_2_2(ch0_coeff_2_2),.coeff_2_3(ch0_coeff_2_3),.coeff_2_4(ch0_coeff_2_4),
	.coeff_2_5(ch0_coeff_2_5),.coeff_2_6(ch0_coeff_2_6),
	.coeff_2_7(ch0_coeff_2_7),.coeff_2_8(ch0_coeff_2_8),.coeff_2_9(ch0_coeff_2_9),.coeff_2_10(ch0_coeff_2_10),
	.coeff_3_0(ch0_coeff_3_0),.coeff_3_1(ch0_coeff_3_1),
	.coeff_3_2(ch0_coeff_3_2),.coeff_3_3(ch0_coeff_3_3),.coeff_3_4(ch0_coeff_3_4),.coeff_3_5(ch0_coeff_3_5),
	.coeff_3_6(ch0_coeff_3_6),.coeff_3_7(ch0_coeff_3_7),
	.coeff_3_8(ch0_coeff_3_8),.coeff_3_9(ch0_coeff_3_9),.coeff_4_0(ch0_coeff_4_0),.coeff_4_1(ch0_coeff_4_1),
	.coeff_4_2(ch0_coeff_4_2),.coeff_4_3(ch0_coeff_4_3),
	.coeff_4_4(ch0_coeff_4_4),.coeff_4_5(ch0_coeff_4_5),.coeff_4_6(ch0_coeff_4_6),.coeff_4_7(ch0_coeff_4_7),
	.coeff_4_8(ch0_coeff_4_8),.coeff_4_9(ch0_coeff_4_9),
	.coeff_4_10(ch0_coeff_4_10),.coeff_3_10(ch0_coeff_3_10),
	.section_select(section_select));	
	
result res (.clk(clk), .reset(reset), .srdyi(srdyo_NLC1ch), .fp_res(fp_res), .srdyo(srdyo), 
            .res_0(ch0_x_lin),
            .res_1(ch1_x_lin),
            .res_2(ch2_x_lin),
            .res_3(ch3_x_lin),
            .res_4(ch4_x_lin),
            .res_5(ch5_x_lin),
            .res_6(ch6_x_lin),
            .res_7(ch7_x_lin),
            .res_8(ch8_x_lin),
            .res_9(ch9_x_lin),
            .res_10(ch10_x_lin),
            .res_11(ch11_x_lin),
            .res_12(ch12_x_lin),
            .res_13(ch13_x_lin),
            .res_14(ch14_x_lin),
            .res_15(ch15_x_lin),
            .res_16(ch16_x_lin),
            .res_17(ch17_x_lin),
            .res_18(ch18_x_lin),
            .res_19(ch19_x_lin),
            .res_20(ch20_x_lin),
            .res_21(ch21_x_lin),
            .res_22(ch22_x_lin),
            .res_23(ch23_x_lin),
            .res_24(ch24_x_lin),
            .res_25(ch25_x_lin),
            .res_26(ch26_x_lin),
            .res_27(ch27_x_lin),
            .res_28(ch28_x_lin),
            .res_29(ch29_x_lin),
            .res_30(ch30_x_lin),
            .res_31(ch31_x_lin)            
);
	

endmodule
